`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:46:30 03/27/2018 
// Design Name: 
// Module Name:    TOP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module TOP(
	input BS_one,
	input BS_zero,
	input PS_top,
	input	Z_top,
	input BrA_top,
	input RAA_top,
	input RC_1_top,
	output MUX_C_out
    );

reg mux_c_select = 
	 
always @(*)
begin
	
end


endmodule
