`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:16:24 03/27/2018 
// Design Name: 
// Module Name:    Mod_Function_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Mod_Function_unit(
	input A,
	input B,
	input SH,
	input FS,
	output Z_out,
	output C_out,
	output N_out,
	output V_out,
	output F
    );


endmodule
